*CTAT Circuit

.lib "../sky130_fd_pr/models/sky130.lib.spice tt"
.include "../sky130_fd_pr/models/sky130_fd_pr__model__pnp.model.spice"


.global vdd gnd
.temp 27

xqp1 gnd gnd qp1 gnd sky130_fd_pr__pnp_05v5_W3p40L3p40

v1 vdd gnd 2
i1 vdd qp1 10u

.dc temp -40 125 5 i1 1.25u 10u 1.25u

.control
run
plot v(qp1)
.endc
.end
